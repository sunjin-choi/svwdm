////==============================================================================
//// Author: Sunjin Choi
//// Description: Virtual Wavelength Probe
//// Signals:
//// Note: 
//// Variable naming conventions:
////    signals => snake_case
////    Parameters (aliasing signal values) => SNAKE_CASE with all caps
////    Parameters (not aliasing signal values) => CamelCase
////==============================================================================
//
//// verilog_format: off
//`timescale 1ns/1ps
//`default_nettype none
//// verilog_format: on
//
//module wprobe #(
//    parameter real Threshold = 0.5
//) (
//
//    // input signals
//    input var waves_t i_phot_waves,
//
//    // output signals
//    output real wavelengths
//);
//
//  // ----------------------------------------------------------------------
//  // Parameters
//  // ----------------------------------------------------------------------
//
//  // ----------------------------------------------------------------------
//
//  // ----------------------------------------------------------------------
//  // Local Parameters
//  // ----------------------------------------------------------------------
//
//  // ----------------------------------------------------------------------
//
//  // ----------------------------------------------------------------------
//  // Inputs / Outputs
//  // ----------------------------------------------------------------------
//
//  // ----------------------------------------------------------------------
//
//  // ----------------------------------------------------------------------
//  // Signals
//  // ----------------------------------------------------------------------
//
//  // ----------------------------------------------------------------------
//
//  // ----------------------------------------------------------------------
//  // Assigns
//  // ----------------------------------------------------------------------
//
//  // ----------------------------------------------------------------------
//
//
//endmodule
//
//`default_nettype wire
//
